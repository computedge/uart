class driver;
	virtual uart_intf.uart_driver vif;

	function new(virtual uart_intf.uart_driver vif);
		this.vif =  vif;
	endfunction



	task reset_signals();
		vif.PSEL 	<= 0;
		vif.PENABLE 	<= 0;
		vif.PWRITE 	<= 0;
		vif.PADDR 	<= 0;
		vif.PWDATA 	<= 0;
	endtask

	task drive (apb_transaction tr);
		@(posedge vif.PCLK)
		vif.PSEL	<= 1;
		vif.PADDR	<= tr.paddr;
		vif.PWRITE	<= tr.write;
		vif.PWDATA	<= tr.pdata;
		vif.PENABLE	<= 0;

		@(posedge vif.PCLK);
		vif.PENABLE	<= 1;
		wait (vif.PREADY);

		@(posedge vif.PCLK);
		vif.PSEL	<= 0;
		vif.PENABLE	<= 0;
		tr.display("DRIVER");
	endtask


  	// Task write
  	task write(string msg = "" , logic [7:0] reg_addr, logic write, logic [7:0] wdata);
  	        tr.message_display(msg);
  	        tr.paddr = reg_addr;
  	        tr.pdata = wdata;
  	        tr.write = write;
  	endtask
endclass
